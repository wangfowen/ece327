library ieee;
use ieee.std_logic_1164.all;

entity add2 is
  port ( i_a, i_b, i_cin : in std_logic;
         o_cout : out std_logic
  );
end add2;

architecture main of add2 is
begin

end architecture;
